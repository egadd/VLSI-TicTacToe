
module ai ( registers, row, col );
  input [17:0] registers;
  output [1:0] row;
  output [1:0] col;
  wire   n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158;

  nor2_1x U86 ( .a(n125), .b(n124), .y(n126) );
  nand2_1x U87 ( .a(n87), .b(n103), .y(n124) );
  nor2_1x U88 ( .a(n109), .b(n84), .y(n127) );
  nor2_1x U89 ( .a(n134), .b(n83), .y(n84) );
  nor2_1x U90 ( .a(n142), .b(n106), .y(n83) );
  nand2_1x U91 ( .a(n138), .b(n120), .y(n121) );
  nor2_1x U92 ( .a(n117), .b(n129), .y(n119) );
  nand2_1x U93 ( .a(n147), .b(n115), .y(n116) );
  inv_1x U94 ( .a(n155), .y(n123) );
  inv_1x U95 ( .a(n152), .y(n154) );
  nand2_1x U96 ( .a(n103), .b(n97), .y(n118) );
  nand2_1x U97 ( .a(n148), .b(n147), .y(n149) );
  nand2_1x U98 ( .a(n143), .b(n142), .y(n144) );
  nor2_1x U99 ( .a(n129), .b(n110), .y(n143) );
  nand2_1x U100 ( .a(n142), .b(n135), .y(n150) );
  nand2_1x U101 ( .a(n136), .b(n134), .y(n151) );
  nor2_1x U102 ( .a(n94), .b(n135), .y(n134) );
  nor2_1x U103 ( .a(n133), .b(n132), .y(n136) );
  inv_1x U104 ( .a(n135), .y(n125) );
  nand2_1x U105 ( .a(n114), .b(n117), .y(n135) );
  inv_4x U106 ( .a(registers[10]), .y(n114) );
  inv_1x U107 ( .a(n153), .y(n112) );
  inv_1x U108 ( .a(n139), .y(n106) );
  inv_1x U109 ( .a(n103), .y(n108) );
  nand2_1x U110 ( .a(n140), .b(n101), .y(n110) );
  inv_1x U111 ( .a(n94), .y(n140) );
  nand2_1x U112 ( .a(n103), .b(n102), .y(n113) );
  nand2_1x U113 ( .a(n97), .b(n96), .y(n98) );
  inv_1x U114 ( .a(n129), .y(n115) );
  nor2_1x U115 ( .a(n94), .b(n141), .y(n97) );
  inv_1x U116 ( .a(n95), .y(n138) );
  inv_1x U117 ( .a(n93), .y(n104) );
  nand2_1x U118 ( .a(n147), .b(n133), .y(n93) );
  inv_1x U119 ( .a(n88), .y(n133) );
  inv_1x U120 ( .a(n87), .y(n147) );
  inv_1x U121 ( .a(n132), .y(n101) );
  nor2_1x U122 ( .a(n109), .b(n142), .y(n103) );
  nor2_2x U123 ( .a(registers[1]), .b(registers[0]), .y(n109) );
  nor2_1x U124 ( .a(registers[10]), .b(n117), .y(n139) );
  nor2_1x U125 ( .a(registers[7]), .b(registers[6]), .y(n129) );
  nor2_1x U126 ( .a(registers[17]), .b(registers[16]), .y(n141) );
  nor2_1x U127 ( .a(registers[3]), .b(registers[2]), .y(n95) );
  nor2_1x U128 ( .a(registers[15]), .b(registers[14]), .y(n88) );
  nor2_1x U129 ( .a(registers[9]), .b(registers[8]), .y(n87) );
  nor2_1x U130 ( .a(registers[5]), .b(registers[4]), .y(n94) );
  nor2_1x U131 ( .a(registers[11]), .b(registers[10]), .y(n132) );
  nor2_1x U132 ( .a(registers[12]), .b(registers[13]), .y(n142) );
  inv_4x U133 ( .a(n109), .y(n158) );
  inv_1x U134 ( .a(registers[13]), .y(n82) );
  a2o1_1x U135 ( .a(registers[6]), .b(n82), .c(registers[12]), .y(n117) );
  nand3_1x U136 ( .a(n127), .b(n101), .c(n93), .y(n92) );
  and2_1x U137 ( .a(n143), .b(n125), .y(n85) );
  a2o1_1x U138 ( .a(n139), .b(n101), .c(n85), .y(n86) );
  nand3_1x U139 ( .a(n103), .b(n95), .c(n86), .y(n91) );
  nand3_1x U140 ( .a(n147), .b(n115), .c(n88), .y(n152) );
  a2o1_1x U141 ( .a(n95), .b(n152), .c(n118), .y(n89) );
  a2o1_1x U142 ( .a(n124), .b(n89), .c(n114), .y(n90) );
  nand3_1x U143 ( .a(n92), .b(n91), .c(n90), .y(col[0]) );
  nand3_1x U144 ( .a(n94), .b(n104), .c(n138), .y(n100) );
  nand3_1x U145 ( .a(n115), .b(n95), .c(n133), .y(n96) );
  nand3_1x U146 ( .a(registers[10]), .b(n147), .c(n98), .y(n99) );
  nand3_1x U147 ( .a(n101), .b(n100), .c(n99), .y(n102) );
  nand3_1x U148 ( .a(n141), .b(n104), .c(n138), .y(n105) );
  a2o1_1x U149 ( .a(n129), .b(n106), .c(n105), .y(n107) );
  nor3_1x U150 ( .a(n110), .b(n108), .c(n107), .y(n153) );
  nand3_1x U151 ( .a(n125), .b(n158), .c(n110), .y(n111) );
  nand3_1x U152 ( .a(n113), .b(n112), .c(n111), .y(col[1]) );
  nor3_1x U153 ( .a(n114), .b(n138), .c(n118), .y(n155) );
  nand3_1x U154 ( .a(n134), .b(n158), .c(n116), .y(n122) );
  nor3_1x U155 ( .a(n119), .b(registers[10]), .c(n118), .y(n120) );
  nand3_1x U156 ( .a(n123), .b(n122), .c(n121), .y(n131) );
  a2o1_1x U157 ( .a(n127), .b(n132), .c(n126), .y(n128) );
  a2o1_1x U158 ( .a(n129), .b(n155), .c(n128), .y(n130) );
  a2o1_1x U159 ( .a(n133), .b(n131), .c(n130), .y(row[0]) );
  or2_1x U160 ( .a(n136), .b(n143), .y(n137) );
  nand3_1x U161 ( .a(n139), .b(n138), .c(n137), .y(n146) );
  nand3_1x U162 ( .a(registers[10]), .b(n141), .c(n140), .y(n145) );
  nand3_1x U163 ( .a(n146), .b(n145), .c(n144), .y(n148) );
  nand3_1x U164 ( .a(n151), .b(n150), .c(n149), .y(n157) );
  a2o1_1x U165 ( .a(n155), .b(n154), .c(n153), .y(n156) );
  a2o1_1x U166 ( .a(n158), .b(n157), .c(n156), .y(row[1]) );
endmodule

