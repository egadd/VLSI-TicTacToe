/home/egadd/VLSI-TicTacToe/verilog/tictactoe.sv