/courses/e158/15/lab3/muddlib.lef